package ast_we_package;

  `include "macro.sv"
  `include "ast_we_transaction.sv"
  `include "ast_we_generator.sv"
  `include "ast_we_driver.sv"
  `include "ast_we_enviroment.sv"

endpackage