package lifo_package;
  `include "defines.svh"
  `include "trans_from_monitor.sv"
  `include "trans_from_generator.sv"
  `include "lifo_generator.sv"
  `include "lifo_driver.sv"
  `include "lifo_monitor.sv"
  `include "lifo_scoreboard.sv"
  `include "lifo_enviroment.sv"
endpackage